magic
tech sky130A
magscale 1 2
timestamp 1658946959
<< obsli1 >>
rect 1104 2159 158884 157777
<< obsm1 >>
rect 106 8 159790 157808
<< metal2 >>
rect 662 159200 718 160000
rect 2042 159200 2098 160000
rect 3422 159200 3478 160000
rect 4802 159200 4858 160000
rect 6274 159200 6330 160000
rect 7654 159200 7710 160000
rect 9034 159200 9090 160000
rect 10414 159200 10470 160000
rect 11886 159200 11942 160000
rect 13266 159200 13322 160000
rect 14646 159200 14702 160000
rect 16026 159200 16082 160000
rect 17498 159200 17554 160000
rect 18878 159200 18934 160000
rect 20258 159200 20314 160000
rect 21638 159200 21694 160000
rect 23110 159200 23166 160000
rect 24490 159200 24546 160000
rect 25870 159200 25926 160000
rect 27250 159200 27306 160000
rect 28722 159200 28778 160000
rect 30102 159200 30158 160000
rect 31482 159200 31538 160000
rect 32862 159200 32918 160000
rect 34334 159200 34390 160000
rect 35714 159200 35770 160000
rect 37094 159200 37150 160000
rect 38474 159200 38530 160000
rect 39946 159200 40002 160000
rect 41326 159200 41382 160000
rect 42706 159200 42762 160000
rect 44086 159200 44142 160000
rect 45558 159200 45614 160000
rect 46938 159200 46994 160000
rect 48318 159200 48374 160000
rect 49698 159200 49754 160000
rect 51170 159200 51226 160000
rect 52550 159200 52606 160000
rect 53930 159200 53986 160000
rect 55310 159200 55366 160000
rect 56782 159200 56838 160000
rect 58162 159200 58218 160000
rect 59542 159200 59598 160000
rect 60922 159200 60978 160000
rect 62394 159200 62450 160000
rect 63774 159200 63830 160000
rect 65154 159200 65210 160000
rect 66534 159200 66590 160000
rect 68006 159200 68062 160000
rect 69386 159200 69442 160000
rect 70766 159200 70822 160000
rect 72146 159200 72202 160000
rect 73618 159200 73674 160000
rect 74998 159200 75054 160000
rect 76378 159200 76434 160000
rect 77758 159200 77814 160000
rect 79230 159200 79286 160000
rect 80610 159200 80666 160000
rect 81990 159200 82046 160000
rect 83462 159200 83518 160000
rect 84842 159200 84898 160000
rect 86222 159200 86278 160000
rect 87602 159200 87658 160000
rect 89074 159200 89130 160000
rect 90454 159200 90510 160000
rect 91834 159200 91890 160000
rect 93214 159200 93270 160000
rect 94686 159200 94742 160000
rect 96066 159200 96122 160000
rect 97446 159200 97502 160000
rect 98826 159200 98882 160000
rect 100298 159200 100354 160000
rect 101678 159200 101734 160000
rect 103058 159200 103114 160000
rect 104438 159200 104494 160000
rect 105910 159200 105966 160000
rect 107290 159200 107346 160000
rect 108670 159200 108726 160000
rect 110050 159200 110106 160000
rect 111522 159200 111578 160000
rect 112902 159200 112958 160000
rect 114282 159200 114338 160000
rect 115662 159200 115718 160000
rect 117134 159200 117190 160000
rect 118514 159200 118570 160000
rect 119894 159200 119950 160000
rect 121274 159200 121330 160000
rect 122746 159200 122802 160000
rect 124126 159200 124182 160000
rect 125506 159200 125562 160000
rect 126886 159200 126942 160000
rect 128358 159200 128414 160000
rect 129738 159200 129794 160000
rect 131118 159200 131174 160000
rect 132498 159200 132554 160000
rect 133970 159200 134026 160000
rect 135350 159200 135406 160000
rect 136730 159200 136786 160000
rect 138110 159200 138166 160000
rect 139582 159200 139638 160000
rect 140962 159200 141018 160000
rect 142342 159200 142398 160000
rect 143722 159200 143778 160000
rect 145194 159200 145250 160000
rect 146574 159200 146630 160000
rect 147954 159200 148010 160000
rect 149334 159200 149390 160000
rect 150806 159200 150862 160000
rect 152186 159200 152242 160000
rect 153566 159200 153622 160000
rect 154946 159200 155002 160000
rect 156418 159200 156474 160000
rect 157798 159200 157854 160000
rect 159178 159200 159234 160000
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2318 0 2374 800
rect 2686 0 2742 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4894 0 4950 800
rect 5262 0 5318 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8206 0 8262 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10414 0 10470 800
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12438 0 12494 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14646 0 14702 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 15934 0 15990 800
rect 16302 0 16358 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17222 0 17278 800
rect 17590 0 17646 800
rect 17958 0 18014 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18878 0 18934 800
rect 19246 0 19302 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20166 0 20222 800
rect 20534 0 20590 800
rect 20810 0 20866 800
rect 21178 0 21234 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24766 0 24822 800
rect 25042 0 25098 800
rect 25410 0 25466 800
rect 25686 0 25742 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 26974 0 27030 800
rect 27342 0 27398 800
rect 27618 0 27674 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28630 0 28686 800
rect 28906 0 28962 800
rect 29274 0 29330 800
rect 29550 0 29606 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30562 0 30618 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32494 0 32550 800
rect 32862 0 32918 800
rect 33138 0 33194 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34150 0 34206 800
rect 34426 0 34482 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35438 0 35494 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36726 0 36782 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37738 0 37794 800
rect 38014 0 38070 800
rect 38382 0 38438 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39670 0 39726 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40590 0 40646 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41602 0 41658 800
rect 41970 0 42026 800
rect 42246 0 42302 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43258 0 43314 800
rect 43534 0 43590 800
rect 43902 0 43958 800
rect 44178 0 44234 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45190 0 45246 800
rect 45466 0 45522 800
rect 45834 0 45890 800
rect 46110 0 46166 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47122 0 47178 800
rect 47398 0 47454 800
rect 47766 0 47822 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49054 0 49110 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50710 0 50766 800
rect 50986 0 51042 800
rect 51354 0 51410 800
rect 51630 0 51686 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52642 0 52698 800
rect 52918 0 52974 800
rect 53286 0 53342 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54942 0 54998 800
rect 55218 0 55274 800
rect 55586 0 55642 800
rect 55862 0 55918 800
rect 56230 0 56286 800
rect 56506 0 56562 800
rect 56874 0 56930 800
rect 57150 0 57206 800
rect 57518 0 57574 800
rect 57794 0 57850 800
rect 58162 0 58218 800
rect 58438 0 58494 800
rect 58806 0 58862 800
rect 59082 0 59138 800
rect 59450 0 59506 800
rect 59818 0 59874 800
rect 60094 0 60150 800
rect 60462 0 60518 800
rect 60738 0 60794 800
rect 61106 0 61162 800
rect 61382 0 61438 800
rect 61750 0 61806 800
rect 62026 0 62082 800
rect 62394 0 62450 800
rect 62670 0 62726 800
rect 63038 0 63094 800
rect 63314 0 63370 800
rect 63682 0 63738 800
rect 63958 0 64014 800
rect 64326 0 64382 800
rect 64602 0 64658 800
rect 64970 0 65026 800
rect 65338 0 65394 800
rect 65614 0 65670 800
rect 65982 0 66038 800
rect 66258 0 66314 800
rect 66626 0 66682 800
rect 66902 0 66958 800
rect 67270 0 67326 800
rect 67546 0 67602 800
rect 67914 0 67970 800
rect 68190 0 68246 800
rect 68558 0 68614 800
rect 68834 0 68890 800
rect 69202 0 69258 800
rect 69478 0 69534 800
rect 69846 0 69902 800
rect 70122 0 70178 800
rect 70490 0 70546 800
rect 70766 0 70822 800
rect 71134 0 71190 800
rect 71502 0 71558 800
rect 71778 0 71834 800
rect 72146 0 72202 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73434 0 73490 800
rect 73710 0 73766 800
rect 74078 0 74134 800
rect 74354 0 74410 800
rect 74722 0 74778 800
rect 74998 0 75054 800
rect 75366 0 75422 800
rect 75642 0 75698 800
rect 76010 0 76066 800
rect 76286 0 76342 800
rect 76654 0 76710 800
rect 76930 0 76986 800
rect 77298 0 77354 800
rect 77666 0 77722 800
rect 77942 0 77998 800
rect 78310 0 78366 800
rect 78586 0 78642 800
rect 78954 0 79010 800
rect 79230 0 79286 800
rect 79598 0 79654 800
rect 79874 0 79930 800
rect 80242 0 80298 800
rect 80518 0 80574 800
rect 80886 0 80942 800
rect 81162 0 81218 800
rect 81530 0 81586 800
rect 81806 0 81862 800
rect 82174 0 82230 800
rect 82450 0 82506 800
rect 82818 0 82874 800
rect 83186 0 83242 800
rect 83462 0 83518 800
rect 83830 0 83886 800
rect 84106 0 84162 800
rect 84474 0 84530 800
rect 84750 0 84806 800
rect 85118 0 85174 800
rect 85394 0 85450 800
rect 85762 0 85818 800
rect 86038 0 86094 800
rect 86406 0 86462 800
rect 86682 0 86738 800
rect 87050 0 87106 800
rect 87326 0 87382 800
rect 87694 0 87750 800
rect 87970 0 88026 800
rect 88338 0 88394 800
rect 88614 0 88670 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89626 0 89682 800
rect 89994 0 90050 800
rect 90270 0 90326 800
rect 90638 0 90694 800
rect 90914 0 90970 800
rect 91282 0 91338 800
rect 91558 0 91614 800
rect 91926 0 91982 800
rect 92202 0 92258 800
rect 92570 0 92626 800
rect 92846 0 92902 800
rect 93214 0 93270 800
rect 93490 0 93546 800
rect 93858 0 93914 800
rect 94134 0 94190 800
rect 94502 0 94558 800
rect 94778 0 94834 800
rect 95146 0 95202 800
rect 95514 0 95570 800
rect 95790 0 95846 800
rect 96158 0 96214 800
rect 96434 0 96490 800
rect 96802 0 96858 800
rect 97078 0 97134 800
rect 97446 0 97502 800
rect 97722 0 97778 800
rect 98090 0 98146 800
rect 98366 0 98422 800
rect 98734 0 98790 800
rect 99010 0 99066 800
rect 99378 0 99434 800
rect 99654 0 99710 800
rect 100022 0 100078 800
rect 100298 0 100354 800
rect 100666 0 100722 800
rect 101034 0 101090 800
rect 101310 0 101366 800
rect 101678 0 101734 800
rect 101954 0 102010 800
rect 102322 0 102378 800
rect 102598 0 102654 800
rect 102966 0 103022 800
rect 103242 0 103298 800
rect 103610 0 103666 800
rect 103886 0 103942 800
rect 104254 0 104310 800
rect 104530 0 104586 800
rect 104898 0 104954 800
rect 105174 0 105230 800
rect 105542 0 105598 800
rect 105818 0 105874 800
rect 106186 0 106242 800
rect 106462 0 106518 800
rect 106830 0 106886 800
rect 107198 0 107254 800
rect 107474 0 107530 800
rect 107842 0 107898 800
rect 108118 0 108174 800
rect 108486 0 108542 800
rect 108762 0 108818 800
rect 109130 0 109186 800
rect 109406 0 109462 800
rect 109774 0 109830 800
rect 110050 0 110106 800
rect 110418 0 110474 800
rect 110694 0 110750 800
rect 111062 0 111118 800
rect 111338 0 111394 800
rect 111706 0 111762 800
rect 111982 0 112038 800
rect 112350 0 112406 800
rect 112718 0 112774 800
rect 112994 0 113050 800
rect 113362 0 113418 800
rect 113638 0 113694 800
rect 114006 0 114062 800
rect 114282 0 114338 800
rect 114650 0 114706 800
rect 114926 0 114982 800
rect 115294 0 115350 800
rect 115570 0 115626 800
rect 115938 0 115994 800
rect 116214 0 116270 800
rect 116582 0 116638 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117502 0 117558 800
rect 117870 0 117926 800
rect 118146 0 118202 800
rect 118514 0 118570 800
rect 118882 0 118938 800
rect 119158 0 119214 800
rect 119526 0 119582 800
rect 119802 0 119858 800
rect 120170 0 120226 800
rect 120446 0 120502 800
rect 120814 0 120870 800
rect 121090 0 121146 800
rect 121458 0 121514 800
rect 121734 0 121790 800
rect 122102 0 122158 800
rect 122378 0 122434 800
rect 122746 0 122802 800
rect 123022 0 123078 800
rect 123390 0 123446 800
rect 123666 0 123722 800
rect 124034 0 124090 800
rect 124310 0 124366 800
rect 124678 0 124734 800
rect 125046 0 125102 800
rect 125322 0 125378 800
rect 125690 0 125746 800
rect 125966 0 126022 800
rect 126334 0 126390 800
rect 126610 0 126666 800
rect 126978 0 127034 800
rect 127254 0 127310 800
rect 127622 0 127678 800
rect 127898 0 127954 800
rect 128266 0 128322 800
rect 128542 0 128598 800
rect 128910 0 128966 800
rect 129186 0 129242 800
rect 129554 0 129610 800
rect 129830 0 129886 800
rect 130198 0 130254 800
rect 130566 0 130622 800
rect 130842 0 130898 800
rect 131210 0 131266 800
rect 131486 0 131542 800
rect 131854 0 131910 800
rect 132130 0 132186 800
rect 132498 0 132554 800
rect 132774 0 132830 800
rect 133142 0 133198 800
rect 133418 0 133474 800
rect 133786 0 133842 800
rect 134062 0 134118 800
rect 134430 0 134486 800
rect 134706 0 134762 800
rect 135074 0 135130 800
rect 135350 0 135406 800
rect 135718 0 135774 800
rect 135994 0 136050 800
rect 136362 0 136418 800
rect 136730 0 136786 800
rect 137006 0 137062 800
rect 137374 0 137430 800
rect 137650 0 137706 800
rect 138018 0 138074 800
rect 138294 0 138350 800
rect 138662 0 138718 800
rect 138938 0 138994 800
rect 139306 0 139362 800
rect 139582 0 139638 800
rect 139950 0 140006 800
rect 140226 0 140282 800
rect 140594 0 140650 800
rect 140870 0 140926 800
rect 141238 0 141294 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142158 0 142214 800
rect 142526 0 142582 800
rect 142894 0 142950 800
rect 143170 0 143226 800
rect 143538 0 143594 800
rect 143814 0 143870 800
rect 144182 0 144238 800
rect 144458 0 144514 800
rect 144826 0 144882 800
rect 145102 0 145158 800
rect 145470 0 145526 800
rect 145746 0 145802 800
rect 146114 0 146170 800
rect 146390 0 146446 800
rect 146758 0 146814 800
rect 147034 0 147090 800
rect 147402 0 147458 800
rect 147678 0 147734 800
rect 148046 0 148102 800
rect 148414 0 148470 800
rect 148690 0 148746 800
rect 149058 0 149114 800
rect 149334 0 149390 800
rect 149702 0 149758 800
rect 149978 0 150034 800
rect 150346 0 150402 800
rect 150622 0 150678 800
rect 150990 0 151046 800
rect 151266 0 151322 800
rect 151634 0 151690 800
rect 151910 0 151966 800
rect 152278 0 152334 800
rect 152554 0 152610 800
rect 152922 0 152978 800
rect 153198 0 153254 800
rect 153566 0 153622 800
rect 153842 0 153898 800
rect 154210 0 154266 800
rect 154578 0 154634 800
rect 154854 0 154910 800
rect 155222 0 155278 800
rect 155498 0 155554 800
rect 155866 0 155922 800
rect 156142 0 156198 800
rect 156510 0 156566 800
rect 156786 0 156842 800
rect 157154 0 157210 800
rect 157430 0 157486 800
rect 157798 0 157854 800
rect 158074 0 158130 800
rect 158442 0 158498 800
rect 158718 0 158774 800
rect 159086 0 159142 800
rect 159362 0 159418 800
rect 159730 0 159786 800
<< obsm2 >>
rect 112 159144 606 159200
rect 774 159144 1986 159200
rect 2154 159144 3366 159200
rect 3534 159144 4746 159200
rect 4914 159144 6218 159200
rect 6386 159144 7598 159200
rect 7766 159144 8978 159200
rect 9146 159144 10358 159200
rect 10526 159144 11830 159200
rect 11998 159144 13210 159200
rect 13378 159144 14590 159200
rect 14758 159144 15970 159200
rect 16138 159144 17442 159200
rect 17610 159144 18822 159200
rect 18990 159144 20202 159200
rect 20370 159144 21582 159200
rect 21750 159144 23054 159200
rect 23222 159144 24434 159200
rect 24602 159144 25814 159200
rect 25982 159144 27194 159200
rect 27362 159144 28666 159200
rect 28834 159144 30046 159200
rect 30214 159144 31426 159200
rect 31594 159144 32806 159200
rect 32974 159144 34278 159200
rect 34446 159144 35658 159200
rect 35826 159144 37038 159200
rect 37206 159144 38418 159200
rect 38586 159144 39890 159200
rect 40058 159144 41270 159200
rect 41438 159144 42650 159200
rect 42818 159144 44030 159200
rect 44198 159144 45502 159200
rect 45670 159144 46882 159200
rect 47050 159144 48262 159200
rect 48430 159144 49642 159200
rect 49810 159144 51114 159200
rect 51282 159144 52494 159200
rect 52662 159144 53874 159200
rect 54042 159144 55254 159200
rect 55422 159144 56726 159200
rect 56894 159144 58106 159200
rect 58274 159144 59486 159200
rect 59654 159144 60866 159200
rect 61034 159144 62338 159200
rect 62506 159144 63718 159200
rect 63886 159144 65098 159200
rect 65266 159144 66478 159200
rect 66646 159144 67950 159200
rect 68118 159144 69330 159200
rect 69498 159144 70710 159200
rect 70878 159144 72090 159200
rect 72258 159144 73562 159200
rect 73730 159144 74942 159200
rect 75110 159144 76322 159200
rect 76490 159144 77702 159200
rect 77870 159144 79174 159200
rect 79342 159144 80554 159200
rect 80722 159144 81934 159200
rect 82102 159144 83406 159200
rect 83574 159144 84786 159200
rect 84954 159144 86166 159200
rect 86334 159144 87546 159200
rect 87714 159144 89018 159200
rect 89186 159144 90398 159200
rect 90566 159144 91778 159200
rect 91946 159144 93158 159200
rect 93326 159144 94630 159200
rect 94798 159144 96010 159200
rect 96178 159144 97390 159200
rect 97558 159144 98770 159200
rect 98938 159144 100242 159200
rect 100410 159144 101622 159200
rect 101790 159144 103002 159200
rect 103170 159144 104382 159200
rect 104550 159144 105854 159200
rect 106022 159144 107234 159200
rect 107402 159144 108614 159200
rect 108782 159144 109994 159200
rect 110162 159144 111466 159200
rect 111634 159144 112846 159200
rect 113014 159144 114226 159200
rect 114394 159144 115606 159200
rect 115774 159144 117078 159200
rect 117246 159144 118458 159200
rect 118626 159144 119838 159200
rect 120006 159144 121218 159200
rect 121386 159144 122690 159200
rect 122858 159144 124070 159200
rect 124238 159144 125450 159200
rect 125618 159144 126830 159200
rect 126998 159144 128302 159200
rect 128470 159144 129682 159200
rect 129850 159144 131062 159200
rect 131230 159144 132442 159200
rect 132610 159144 133914 159200
rect 134082 159144 135294 159200
rect 135462 159144 136674 159200
rect 136842 159144 138054 159200
rect 138222 159144 139526 159200
rect 139694 159144 140906 159200
rect 141074 159144 142286 159200
rect 142454 159144 143666 159200
rect 143834 159144 145138 159200
rect 145306 159144 146518 159200
rect 146686 159144 147898 159200
rect 148066 159144 149278 159200
rect 149446 159144 150750 159200
rect 150918 159144 152130 159200
rect 152298 159144 153510 159200
rect 153678 159144 154890 159200
rect 155058 159144 156362 159200
rect 156530 159144 157742 159200
rect 157910 159144 159122 159200
rect 159290 159144 159784 159200
rect 112 856 159784 159144
rect 222 2 330 856
rect 498 2 698 856
rect 866 2 974 856
rect 1142 2 1342 856
rect 1510 2 1618 856
rect 1786 2 1986 856
rect 2154 2 2262 856
rect 2430 2 2630 856
rect 2798 2 2906 856
rect 3074 2 3274 856
rect 3442 2 3550 856
rect 3718 2 3918 856
rect 4086 2 4194 856
rect 4362 2 4562 856
rect 4730 2 4838 856
rect 5006 2 5206 856
rect 5374 2 5482 856
rect 5650 2 5850 856
rect 6018 2 6218 856
rect 6386 2 6494 856
rect 6662 2 6862 856
rect 7030 2 7138 856
rect 7306 2 7506 856
rect 7674 2 7782 856
rect 7950 2 8150 856
rect 8318 2 8426 856
rect 8594 2 8794 856
rect 8962 2 9070 856
rect 9238 2 9438 856
rect 9606 2 9714 856
rect 9882 2 10082 856
rect 10250 2 10358 856
rect 10526 2 10726 856
rect 10894 2 11002 856
rect 11170 2 11370 856
rect 11538 2 11646 856
rect 11814 2 12014 856
rect 12182 2 12382 856
rect 12550 2 12658 856
rect 12826 2 13026 856
rect 13194 2 13302 856
rect 13470 2 13670 856
rect 13838 2 13946 856
rect 14114 2 14314 856
rect 14482 2 14590 856
rect 14758 2 14958 856
rect 15126 2 15234 856
rect 15402 2 15602 856
rect 15770 2 15878 856
rect 16046 2 16246 856
rect 16414 2 16522 856
rect 16690 2 16890 856
rect 17058 2 17166 856
rect 17334 2 17534 856
rect 17702 2 17902 856
rect 18070 2 18178 856
rect 18346 2 18546 856
rect 18714 2 18822 856
rect 18990 2 19190 856
rect 19358 2 19466 856
rect 19634 2 19834 856
rect 20002 2 20110 856
rect 20278 2 20478 856
rect 20646 2 20754 856
rect 20922 2 21122 856
rect 21290 2 21398 856
rect 21566 2 21766 856
rect 21934 2 22042 856
rect 22210 2 22410 856
rect 22578 2 22686 856
rect 22854 2 23054 856
rect 23222 2 23330 856
rect 23498 2 23698 856
rect 23866 2 24066 856
rect 24234 2 24342 856
rect 24510 2 24710 856
rect 24878 2 24986 856
rect 25154 2 25354 856
rect 25522 2 25630 856
rect 25798 2 25998 856
rect 26166 2 26274 856
rect 26442 2 26642 856
rect 26810 2 26918 856
rect 27086 2 27286 856
rect 27454 2 27562 856
rect 27730 2 27930 856
rect 28098 2 28206 856
rect 28374 2 28574 856
rect 28742 2 28850 856
rect 29018 2 29218 856
rect 29386 2 29494 856
rect 29662 2 29862 856
rect 30030 2 30230 856
rect 30398 2 30506 856
rect 30674 2 30874 856
rect 31042 2 31150 856
rect 31318 2 31518 856
rect 31686 2 31794 856
rect 31962 2 32162 856
rect 32330 2 32438 856
rect 32606 2 32806 856
rect 32974 2 33082 856
rect 33250 2 33450 856
rect 33618 2 33726 856
rect 33894 2 34094 856
rect 34262 2 34370 856
rect 34538 2 34738 856
rect 34906 2 35014 856
rect 35182 2 35382 856
rect 35550 2 35750 856
rect 35918 2 36026 856
rect 36194 2 36394 856
rect 36562 2 36670 856
rect 36838 2 37038 856
rect 37206 2 37314 856
rect 37482 2 37682 856
rect 37850 2 37958 856
rect 38126 2 38326 856
rect 38494 2 38602 856
rect 38770 2 38970 856
rect 39138 2 39246 856
rect 39414 2 39614 856
rect 39782 2 39890 856
rect 40058 2 40258 856
rect 40426 2 40534 856
rect 40702 2 40902 856
rect 41070 2 41178 856
rect 41346 2 41546 856
rect 41714 2 41914 856
rect 42082 2 42190 856
rect 42358 2 42558 856
rect 42726 2 42834 856
rect 43002 2 43202 856
rect 43370 2 43478 856
rect 43646 2 43846 856
rect 44014 2 44122 856
rect 44290 2 44490 856
rect 44658 2 44766 856
rect 44934 2 45134 856
rect 45302 2 45410 856
rect 45578 2 45778 856
rect 45946 2 46054 856
rect 46222 2 46422 856
rect 46590 2 46698 856
rect 46866 2 47066 856
rect 47234 2 47342 856
rect 47510 2 47710 856
rect 47878 2 48078 856
rect 48246 2 48354 856
rect 48522 2 48722 856
rect 48890 2 48998 856
rect 49166 2 49366 856
rect 49534 2 49642 856
rect 49810 2 50010 856
rect 50178 2 50286 856
rect 50454 2 50654 856
rect 50822 2 50930 856
rect 51098 2 51298 856
rect 51466 2 51574 856
rect 51742 2 51942 856
rect 52110 2 52218 856
rect 52386 2 52586 856
rect 52754 2 52862 856
rect 53030 2 53230 856
rect 53398 2 53598 856
rect 53766 2 53874 856
rect 54042 2 54242 856
rect 54410 2 54518 856
rect 54686 2 54886 856
rect 55054 2 55162 856
rect 55330 2 55530 856
rect 55698 2 55806 856
rect 55974 2 56174 856
rect 56342 2 56450 856
rect 56618 2 56818 856
rect 56986 2 57094 856
rect 57262 2 57462 856
rect 57630 2 57738 856
rect 57906 2 58106 856
rect 58274 2 58382 856
rect 58550 2 58750 856
rect 58918 2 59026 856
rect 59194 2 59394 856
rect 59562 2 59762 856
rect 59930 2 60038 856
rect 60206 2 60406 856
rect 60574 2 60682 856
rect 60850 2 61050 856
rect 61218 2 61326 856
rect 61494 2 61694 856
rect 61862 2 61970 856
rect 62138 2 62338 856
rect 62506 2 62614 856
rect 62782 2 62982 856
rect 63150 2 63258 856
rect 63426 2 63626 856
rect 63794 2 63902 856
rect 64070 2 64270 856
rect 64438 2 64546 856
rect 64714 2 64914 856
rect 65082 2 65282 856
rect 65450 2 65558 856
rect 65726 2 65926 856
rect 66094 2 66202 856
rect 66370 2 66570 856
rect 66738 2 66846 856
rect 67014 2 67214 856
rect 67382 2 67490 856
rect 67658 2 67858 856
rect 68026 2 68134 856
rect 68302 2 68502 856
rect 68670 2 68778 856
rect 68946 2 69146 856
rect 69314 2 69422 856
rect 69590 2 69790 856
rect 69958 2 70066 856
rect 70234 2 70434 856
rect 70602 2 70710 856
rect 70878 2 71078 856
rect 71246 2 71446 856
rect 71614 2 71722 856
rect 71890 2 72090 856
rect 72258 2 72366 856
rect 72534 2 72734 856
rect 72902 2 73010 856
rect 73178 2 73378 856
rect 73546 2 73654 856
rect 73822 2 74022 856
rect 74190 2 74298 856
rect 74466 2 74666 856
rect 74834 2 74942 856
rect 75110 2 75310 856
rect 75478 2 75586 856
rect 75754 2 75954 856
rect 76122 2 76230 856
rect 76398 2 76598 856
rect 76766 2 76874 856
rect 77042 2 77242 856
rect 77410 2 77610 856
rect 77778 2 77886 856
rect 78054 2 78254 856
rect 78422 2 78530 856
rect 78698 2 78898 856
rect 79066 2 79174 856
rect 79342 2 79542 856
rect 79710 2 79818 856
rect 79986 2 80186 856
rect 80354 2 80462 856
rect 80630 2 80830 856
rect 80998 2 81106 856
rect 81274 2 81474 856
rect 81642 2 81750 856
rect 81918 2 82118 856
rect 82286 2 82394 856
rect 82562 2 82762 856
rect 82930 2 83130 856
rect 83298 2 83406 856
rect 83574 2 83774 856
rect 83942 2 84050 856
rect 84218 2 84418 856
rect 84586 2 84694 856
rect 84862 2 85062 856
rect 85230 2 85338 856
rect 85506 2 85706 856
rect 85874 2 85982 856
rect 86150 2 86350 856
rect 86518 2 86626 856
rect 86794 2 86994 856
rect 87162 2 87270 856
rect 87438 2 87638 856
rect 87806 2 87914 856
rect 88082 2 88282 856
rect 88450 2 88558 856
rect 88726 2 88926 856
rect 89094 2 89294 856
rect 89462 2 89570 856
rect 89738 2 89938 856
rect 90106 2 90214 856
rect 90382 2 90582 856
rect 90750 2 90858 856
rect 91026 2 91226 856
rect 91394 2 91502 856
rect 91670 2 91870 856
rect 92038 2 92146 856
rect 92314 2 92514 856
rect 92682 2 92790 856
rect 92958 2 93158 856
rect 93326 2 93434 856
rect 93602 2 93802 856
rect 93970 2 94078 856
rect 94246 2 94446 856
rect 94614 2 94722 856
rect 94890 2 95090 856
rect 95258 2 95458 856
rect 95626 2 95734 856
rect 95902 2 96102 856
rect 96270 2 96378 856
rect 96546 2 96746 856
rect 96914 2 97022 856
rect 97190 2 97390 856
rect 97558 2 97666 856
rect 97834 2 98034 856
rect 98202 2 98310 856
rect 98478 2 98678 856
rect 98846 2 98954 856
rect 99122 2 99322 856
rect 99490 2 99598 856
rect 99766 2 99966 856
rect 100134 2 100242 856
rect 100410 2 100610 856
rect 100778 2 100978 856
rect 101146 2 101254 856
rect 101422 2 101622 856
rect 101790 2 101898 856
rect 102066 2 102266 856
rect 102434 2 102542 856
rect 102710 2 102910 856
rect 103078 2 103186 856
rect 103354 2 103554 856
rect 103722 2 103830 856
rect 103998 2 104198 856
rect 104366 2 104474 856
rect 104642 2 104842 856
rect 105010 2 105118 856
rect 105286 2 105486 856
rect 105654 2 105762 856
rect 105930 2 106130 856
rect 106298 2 106406 856
rect 106574 2 106774 856
rect 106942 2 107142 856
rect 107310 2 107418 856
rect 107586 2 107786 856
rect 107954 2 108062 856
rect 108230 2 108430 856
rect 108598 2 108706 856
rect 108874 2 109074 856
rect 109242 2 109350 856
rect 109518 2 109718 856
rect 109886 2 109994 856
rect 110162 2 110362 856
rect 110530 2 110638 856
rect 110806 2 111006 856
rect 111174 2 111282 856
rect 111450 2 111650 856
rect 111818 2 111926 856
rect 112094 2 112294 856
rect 112462 2 112662 856
rect 112830 2 112938 856
rect 113106 2 113306 856
rect 113474 2 113582 856
rect 113750 2 113950 856
rect 114118 2 114226 856
rect 114394 2 114594 856
rect 114762 2 114870 856
rect 115038 2 115238 856
rect 115406 2 115514 856
rect 115682 2 115882 856
rect 116050 2 116158 856
rect 116326 2 116526 856
rect 116694 2 116802 856
rect 116970 2 117170 856
rect 117338 2 117446 856
rect 117614 2 117814 856
rect 117982 2 118090 856
rect 118258 2 118458 856
rect 118626 2 118826 856
rect 118994 2 119102 856
rect 119270 2 119470 856
rect 119638 2 119746 856
rect 119914 2 120114 856
rect 120282 2 120390 856
rect 120558 2 120758 856
rect 120926 2 121034 856
rect 121202 2 121402 856
rect 121570 2 121678 856
rect 121846 2 122046 856
rect 122214 2 122322 856
rect 122490 2 122690 856
rect 122858 2 122966 856
rect 123134 2 123334 856
rect 123502 2 123610 856
rect 123778 2 123978 856
rect 124146 2 124254 856
rect 124422 2 124622 856
rect 124790 2 124990 856
rect 125158 2 125266 856
rect 125434 2 125634 856
rect 125802 2 125910 856
rect 126078 2 126278 856
rect 126446 2 126554 856
rect 126722 2 126922 856
rect 127090 2 127198 856
rect 127366 2 127566 856
rect 127734 2 127842 856
rect 128010 2 128210 856
rect 128378 2 128486 856
rect 128654 2 128854 856
rect 129022 2 129130 856
rect 129298 2 129498 856
rect 129666 2 129774 856
rect 129942 2 130142 856
rect 130310 2 130510 856
rect 130678 2 130786 856
rect 130954 2 131154 856
rect 131322 2 131430 856
rect 131598 2 131798 856
rect 131966 2 132074 856
rect 132242 2 132442 856
rect 132610 2 132718 856
rect 132886 2 133086 856
rect 133254 2 133362 856
rect 133530 2 133730 856
rect 133898 2 134006 856
rect 134174 2 134374 856
rect 134542 2 134650 856
rect 134818 2 135018 856
rect 135186 2 135294 856
rect 135462 2 135662 856
rect 135830 2 135938 856
rect 136106 2 136306 856
rect 136474 2 136674 856
rect 136842 2 136950 856
rect 137118 2 137318 856
rect 137486 2 137594 856
rect 137762 2 137962 856
rect 138130 2 138238 856
rect 138406 2 138606 856
rect 138774 2 138882 856
rect 139050 2 139250 856
rect 139418 2 139526 856
rect 139694 2 139894 856
rect 140062 2 140170 856
rect 140338 2 140538 856
rect 140706 2 140814 856
rect 140982 2 141182 856
rect 141350 2 141458 856
rect 141626 2 141826 856
rect 141994 2 142102 856
rect 142270 2 142470 856
rect 142638 2 142838 856
rect 143006 2 143114 856
rect 143282 2 143482 856
rect 143650 2 143758 856
rect 143926 2 144126 856
rect 144294 2 144402 856
rect 144570 2 144770 856
rect 144938 2 145046 856
rect 145214 2 145414 856
rect 145582 2 145690 856
rect 145858 2 146058 856
rect 146226 2 146334 856
rect 146502 2 146702 856
rect 146870 2 146978 856
rect 147146 2 147346 856
rect 147514 2 147622 856
rect 147790 2 147990 856
rect 148158 2 148358 856
rect 148526 2 148634 856
rect 148802 2 149002 856
rect 149170 2 149278 856
rect 149446 2 149646 856
rect 149814 2 149922 856
rect 150090 2 150290 856
rect 150458 2 150566 856
rect 150734 2 150934 856
rect 151102 2 151210 856
rect 151378 2 151578 856
rect 151746 2 151854 856
rect 152022 2 152222 856
rect 152390 2 152498 856
rect 152666 2 152866 856
rect 153034 2 153142 856
rect 153310 2 153510 856
rect 153678 2 153786 856
rect 153954 2 154154 856
rect 154322 2 154522 856
rect 154690 2 154798 856
rect 154966 2 155166 856
rect 155334 2 155442 856
rect 155610 2 155810 856
rect 155978 2 156086 856
rect 156254 2 156454 856
rect 156622 2 156730 856
rect 156898 2 157098 856
rect 157266 2 157374 856
rect 157542 2 157742 856
rect 157910 2 158018 856
rect 158186 2 158386 856
rect 158554 2 158662 856
rect 158830 2 159030 856
rect 159198 2 159306 856
rect 159474 2 159674 856
<< metal3 >>
rect 159200 79976 160000 80096
<< obsm3 >>
rect 1485 1395 158128 157793
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
rect 111728 2128 112048 157808
rect 127088 2128 127408 157808
rect 142448 2128 142768 157808
rect 157808 2128 158128 157808
<< obsm4 >>
rect 4659 2048 19488 145077
rect 19968 2048 34848 145077
rect 35328 2048 50208 145077
rect 50688 2048 65568 145077
rect 66048 2048 80928 145077
rect 81408 2048 96288 145077
rect 96768 2048 111648 145077
rect 112128 2048 127008 145077
rect 127488 2048 142368 145077
rect 142848 2048 143829 145077
rect 4659 1667 143829 2048
<< labels >>
rlabel metal2 s 662 159200 718 160000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 42706 159200 42762 160000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 46938 159200 46994 160000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 51170 159200 51226 160000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 55310 159200 55366 160000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 59542 159200 59598 160000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 63774 159200 63830 160000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 68006 159200 68062 160000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 72146 159200 72202 160000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 76378 159200 76434 160000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 80610 159200 80666 160000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 4802 159200 4858 160000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 84842 159200 84898 160000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 89074 159200 89130 160000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 93214 159200 93270 160000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 97446 159200 97502 160000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 101678 159200 101734 160000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 105910 159200 105966 160000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 110050 159200 110106 160000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 114282 159200 114338 160000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 118514 159200 118570 160000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 122746 159200 122802 160000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 9034 159200 9090 160000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 126886 159200 126942 160000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 131118 159200 131174 160000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 135350 159200 135406 160000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 139582 159200 139638 160000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 143722 159200 143778 160000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 147954 159200 148010 160000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 152186 159200 152242 160000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 156418 159200 156474 160000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 13266 159200 13322 160000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 17498 159200 17554 160000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 21638 159200 21694 160000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 25870 159200 25926 160000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 30102 159200 30158 160000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 34334 159200 34390 160000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 38474 159200 38530 160000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2042 159200 2098 160000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 44086 159200 44142 160000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 48318 159200 48374 160000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 52550 159200 52606 160000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 56782 159200 56838 160000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 60922 159200 60978 160000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 65154 159200 65210 160000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 69386 159200 69442 160000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 73618 159200 73674 160000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 77758 159200 77814 160000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 81990 159200 82046 160000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 6274 159200 6330 160000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 86222 159200 86278 160000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 90454 159200 90510 160000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 94686 159200 94742 160000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 98826 159200 98882 160000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 103058 159200 103114 160000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 107290 159200 107346 160000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 111522 159200 111578 160000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 115662 159200 115718 160000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 119894 159200 119950 160000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 124126 159200 124182 160000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 10414 159200 10470 160000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 128358 159200 128414 160000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 132498 159200 132554 160000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 136730 159200 136786 160000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 140962 159200 141018 160000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 145194 159200 145250 160000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 149334 159200 149390 160000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 153566 159200 153622 160000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 157798 159200 157854 160000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 14646 159200 14702 160000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 18878 159200 18934 160000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 23110 159200 23166 160000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 27250 159200 27306 160000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 31482 159200 31538 160000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 35714 159200 35770 160000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 39946 159200 40002 160000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3422 159200 3478 160000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 45558 159200 45614 160000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 49698 159200 49754 160000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 53930 159200 53986 160000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 58162 159200 58218 160000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 62394 159200 62450 160000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 66534 159200 66590 160000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 70766 159200 70822 160000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 74998 159200 75054 160000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 79230 159200 79286 160000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 83462 159200 83518 160000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 7654 159200 7710 160000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 87602 159200 87658 160000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 91834 159200 91890 160000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 96066 159200 96122 160000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 100298 159200 100354 160000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 104438 159200 104494 160000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 108670 159200 108726 160000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 112902 159200 112958 160000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 117134 159200 117190 160000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 121274 159200 121330 160000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 125506 159200 125562 160000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 11886 159200 11942 160000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 129738 159200 129794 160000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 133970 159200 134026 160000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 138110 159200 138166 160000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 142342 159200 142398 160000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 146574 159200 146630 160000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 150806 159200 150862 160000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 154946 159200 155002 160000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 159178 159200 159234 160000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 16026 159200 16082 160000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 20258 159200 20314 160000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 24490 159200 24546 160000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 28722 159200 28778 160000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 32862 159200 32918 160000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 37094 159200 37150 160000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 41326 159200 41382 160000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 159362 0 159418 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 159730 0 159786 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 147402 0 147458 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 148414 0 148470 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 149334 0 149390 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 150346 0 150402 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 105542 0 105598 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 124034 0 124090 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 133142 0 133198 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 134062 0 134118 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 135074 0 135130 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 135994 0 136050 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 137006 0 137062 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 138018 0 138074 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 138938 0 138994 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 140870 0 140926 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 143814 0 143870 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 145746 0 145802 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 146758 0 146814 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 147678 0 147734 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 148690 0 148746 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 149702 0 149758 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 150622 0 150678 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 151634 0 151690 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 152554 0 152610 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 153566 0 153622 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 154578 0 154634 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 155498 0 155554 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 78586 0 78642 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 83462 0 83518 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 88338 0 88394 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 90270 0 90326 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 94134 0 94190 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 96158 0 96214 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 97078 0 97134 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 100022 0 100078 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 101954 0 102010 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 121458 0 121514 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 122378 0 122434 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 123390 0 123446 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 124310 0 124366 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 126334 0 126390 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 129186 0 129242 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 134430 0 134486 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 140226 0 140282 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 146114 0 146170 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 129554 0 129610 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal3 s 159200 79976 160000 80096 6 user_clock2
port 502 nsew signal input
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 503 nsew power input
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 503 nsew power input
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 503 nsew power input
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 503 nsew power input
rlabel metal4 s 127088 2128 127408 157808 6 vccd1
port 503 nsew power input
rlabel metal4 s 157808 2128 158128 157808 6 vccd1
port 503 nsew power input
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 504 nsew ground input
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 504 nsew ground input
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 504 nsew ground input
rlabel metal4 s 111728 2128 112048 157808 6 vssd1
port 504 nsew ground input
rlabel metal4 s 142448 2128 142768 157808 6 vssd1
port 504 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 505 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 506 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_ack_o
port 507 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 wbs_adr_i[0]
port 508 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[10]
port 509 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[11]
port 510 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_adr_i[12]
port 511 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_adr_i[13]
port 512 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_adr_i[14]
port 513 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[15]
port 514 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_adr_i[16]
port 515 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_adr_i[17]
port 516 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 wbs_adr_i[18]
port 517 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_adr_i[19]
port 518 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_adr_i[1]
port 519 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_adr_i[20]
port 520 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[21]
port 521 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_adr_i[22]
port 522 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_adr_i[23]
port 523 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_adr_i[24]
port 524 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wbs_adr_i[25]
port 525 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[26]
port 526 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[27]
port 527 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_adr_i[28]
port 528 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_adr_i[29]
port 529 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_adr_i[2]
port 530 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_adr_i[30]
port 531 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_adr_i[31]
port 532 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_adr_i[3]
port 533 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_adr_i[4]
port 534 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[5]
port 535 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[6]
port 536 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_adr_i[7]
port 537 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_adr_i[8]
port 538 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_adr_i[9]
port 539 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_cyc_i
port 540 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_dat_i[0]
port 541 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_i[10]
port 542 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_i[11]
port 543 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_i[12]
port 544 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_i[13]
port 545 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_i[14]
port 546 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_i[15]
port 547 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[16]
port 548 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_i[17]
port 549 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_i[18]
port 550 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_i[19]
port 551 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_i[1]
port 552 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_i[20]
port 553 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_i[21]
port 554 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_i[22]
port 555 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[23]
port 556 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_i[24]
port 557 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_i[25]
port 558 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_i[26]
port 559 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[27]
port 560 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_i[28]
port 561 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_i[29]
port 562 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_i[2]
port 563 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_i[30]
port 564 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_i[31]
port 565 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_i[3]
port 566 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_i[4]
port 567 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[5]
port 568 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[6]
port 569 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_i[7]
port 570 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[8]
port 571 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_i[9]
port 572 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_o[0]
port 573 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_o[10]
port 574 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_o[11]
port 575 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_o[12]
port 576 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_o[13]
port 577 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_o[14]
port 578 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_o[15]
port 579 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[16]
port 580 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_o[17]
port 581 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_o[18]
port 582 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_o[19]
port 583 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 wbs_dat_o[1]
port 584 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[20]
port 585 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_o[21]
port 586 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[22]
port 587 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_o[23]
port 588 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_o[24]
port 589 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 wbs_dat_o[25]
port 590 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_o[26]
port 591 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[27]
port 592 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_o[28]
port 593 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[29]
port 594 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_o[2]
port 595 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_o[30]
port 596 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 wbs_dat_o[31]
port 597 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[3]
port 598 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_o[4]
port 599 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[5]
port 600 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[6]
port 601 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[7]
port 602 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[8]
port 603 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_o[9]
port 604 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 wbs_sel_i[0]
port 605 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_sel_i[1]
port 606 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_sel_i[2]
port 607 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_sel_i[3]
port 608 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_stb_i
port 609 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_we_i
port 610 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 160000 160000
string LEFview TRUE
string GDS_FILE /home/shuttle/space_controller/openlane/user_proj_example/runs/user_proj_example/results/finishing/user_proj_example.gds
string GDS_END 57013094
string GDS_START 834868
<< end >>

